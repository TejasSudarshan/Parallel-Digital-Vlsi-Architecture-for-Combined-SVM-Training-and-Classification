010001110
00000000-1
010101011
00000000-1
010111010
000000001
011000011
000000001
011000111
000000001
010001111
00000000-1
101010101
000000001
001001111
00000000-1
001011001
00000000-1
011101101
000000001
011011001
000000001
010101001
000000001
001100100
000000001
011000111
000000001
010011011
00000000-1
010010001
00000000-1
010111000
000000001
011000001
000000001
101000100
000000001
101001101
000000001
001010111
00000000-1
001111011
00000000-1
101000001
000000001
110011100
000000001
110011001
000000001
111111001
000000001
100011111
000000001
101001100
000000001
000110101
00000000-1
100101010
000000001
011011110
000000001
010110010
00000000-1
100011011
000000001
011010100
000000001
011110011
000000001
001101111
00000000-1
001110001
00000000-1
010010100
00000000-1
001101111
00000000-1
001100101
00000000-1
001100111
00000000-1
001100011
00000000-1
011001000
000000001
001001100
00000000-1
001111011
00000000-1
010000100
00000000-1
001010111
00000000-1
011001001
000000001
000111000
00000000-1
011010011
000000001
